entity test is
   port (i0, i1 : in bit; ci : in bit; s : out bit; co : out bit);
 end test;
 
 architecture rtl of test is
 begin
 end rtl;