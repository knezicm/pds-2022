
`ifndef __FOUR_BIT_FULL_ADDER_DEFINES_SVH__
`define __FOUR_BIT_FULL_ADDER_DEFINES_SVH__

`ifndef FBDA_X_WIDTH
    `define FBDA_X_WIDTH 4
`endif /* FBDA_X_WIDTH */

`ifndef FBDA_Y_WIDTH
    `define FBDA_Y_WIDTH 4
`endif /* FBDA_Y_WIDTH */

`ifndef FBDA_RES_WIDTH
    `define FBDA_RES_WIDTH 4
`endif /* FBDA_RES_WIDTH */

`ifndef FBDA_C_WIDTH
    `define FBDA_C_WIDTH 2
    `define FBDA_C_IN    0
    `define FBDA_C_OUT   1
`endif /* FBDA_C_WIDTH */


`endif /* __FOUR_BIT_FULL_ADDER_DEFINES_SVH__ */
