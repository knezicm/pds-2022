library ieee;
use ieee.std_logic_1164.all;

entity prio_encoder is
	port(
		r : in std_logic_vector(3 downto 0);
		code : out std_logic_vector(1 downto 0);
		active : out std_logic
	);
end prio_encoder;

architecture cond_arch of prio_encoder is
begin
	code <=	"11" when (r(3) = '1') else
				"10" when (r(2) = '1') else
				"01" when (r(1) = '1') else
				"00";
	
	active <= r(3) or r(2) or r(1) or r(0);
end cond_arch;

architecture sel_arch of prio_encoder is
begin
	with r select
		code <=	"11" 	when 	"1000"|"1001"|"1010"|"1011"|
									"1100"|"1101"|"1110"|"1111",
					"10" 	when	"0100"|"0101"|"0110"|"0111",
					"01" 	when	"0010"|"0011",
					"00"	when	others;
	
	active <= r(3) or r(2) or r(1) or r(0);
end sel_arch;

configuration prio_encoder_cfg of prio_encoder is
	for sel_arch
	end for;
end prio_encoder_cfg;
