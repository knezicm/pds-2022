library ieee;
use ieee.std_logic_1164.all;

entity test is


	port
	(
		
		x	: in  std_logic_vector(7 downto 0);
		
		y	: out std_logic
		
	);
end test;


architecture test_arch of test is

begin

	

end test_arch;
