
`ifndef __FOUR_BIT_FULL_SUBTRACTOR_DEFINES_SVH__
`define __FOUR_BIT_FULL_SUBTRACTOR_DEFINES_SVH__

`ifndef FBFS_X_WIDTH
    `define FBFS_X_WIDTH 4
`endif /* FBFS_X_WIDTH */

`ifndef FBFS_Y_WIDTH
    `define FBFS_Y_WIDTH 4
`endif /* FBFS_Y_WIDTH */

`ifndef FBFS_D_WIDTH
    `define FBFS_D_WIDTH 4
`endif /* FBFS_D_WIDTH */

`ifndef FBFS_B_WIDTH
    `define FBFS_B_WIDTH 2
    `define FBFS_B_IN    0
    `define FBFS_B_OUT   1
`endif /* FBFS_B_WIDTH*/


`endif /* __FOUR_BIT_FULL_SUBTRACTOR_DEFINES_SVH__ */
