library ieee;
use ieee.std_logic_1164.all;


entity test is
port (

	input  : in std_logic_vector (3 downto 0);
	sel    : in std_logic_vector (1 downto 0);
	output : out std_logic
	);
end test;

architecture test_arch of test is
	
end test_arch;
