
`ifndef __NAND2_DEFINES_SVH__
`define __NAND2_DEFINES_SVH__

`ifndef NAND2_IN_WIDTH
    `define NAND2_IN_WIDTH          2
    `define NAND2_A                 0
    `define NAND2_B                 1
`endif /* NAND2_IN_WIDTH */

`ifndef NAND2_OUT_WIDTH
    `define NAND2_OUT_WIDTH         1
    `define NAND2_Y                 0   
`endif /* NAND2_OUT_WIDTH */

`endif /* __NAND2_DEFINES_SVH__ */
