library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity simple_alu is
	port(
		ctrl : in std_logic_vector(2 downto 0);
		src0, src1 : in std_logic_vector(7 downto 0);
		result : out std_logic_vector(7 downto 0)
	);
end simple_alu;

architecture cond_arch of simple_alu is
	signal sum, diff, inc : std_logic_vector(7 downto 0);
begin
	sum <= std_logic_vector(signed(src0) + signed(src1));
	diff <= std_logic_vector(signed(src0) - signed(src1));
	inc <= std_logic_vector(signed(src0) + 1);
	
	result <= 	inc	when ctrl(2) = '0' else
					sum	when ctrl(1 downto 0) = "00" else
					diff	when ctrl(1 downto 0) = "01" else
					src0 and src1 when ctrl(1 downto 0) = "10" else
					src0 or src1;
end cond_arch;

architecture sel_arch of simple_alu is
	signal sum, diff, inc : std_logic_vector(7 downto 0);
begin
	sum <= std_logic_vector(signed(src0) + signed(src1));
	diff <= std_logic_vector(signed(src0) - signed(src1));
	inc <= std_logic_vector(signed(src0) + 1);
	
	with ctrl select
		result <= 	inc				when "000"|"001"|"010"|"011",
						sum				when "100",
						diff				when "101",
						src0 and src1	when "110",
						src0 or src1	when others;	-- "111"
end sel_arch;

configuration simple_alu_cfg of simple_alu is
	for sel_arch
	end for;
end simple_alu_cfg;
