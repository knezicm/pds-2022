  -----------------------------------------------------------------------------
  -- Faculty of Electrical Engineering
  -- PDS 2022
  -- https://github.com/knezicm/pds-2022/
  -----------------------------------------------------------------------------
  --
  -- unit name:     NAND2
  --
  -- description:
  --
  --   This file implements a simple NAND2 logic.
  --
  -----------------------------------------------------------------------------
  -- Copyright (c) 2022 Faculty of Electrical Engineering
  -----------------------------------------------------------------------------
  -- The MIT License
  -----------------------------------------------------------------------------
  -- Copyright 2022 Faculty of Electrical Engineering
  --
  -- Permission is hereby granted, free of charge, to any person obtaining a
  -- copy of this software and associated documentation files (the "Software"),
  -- to deal in the Software without restriction, including without limitation
  -- the rights to use, copy, modify, merge, publish, distribute, sublicense,
  -- and/or sell copies of the Software, and to permit persons to whom
  -- the Software is furnished to do so, subject to the following conditions:
  --
  -- The above copyright notice and this permission notice shall be included in
  -- all copies or substantial portions of the Software.
  --
  -- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
  -- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
  -- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
  -- THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
  -- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
  -- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
  -- OTHER DEALINGS IN THE SOFTWARE
  -----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity nand2 is
port (
  A_i : in  std_logic;
  B_i : in  std_logic;
  Y_o : out std_logic
);
end nand2;

architecture arch of nand2 is
begin
  Y_o <= A_i nand B_i;
end behav;
